* Equivalent circuit model for E:\touchstone_files\vccline.ckt
.SUBCKT vccline po1 po2
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Vsp2 po2 p2 0
Vsr2 p2 pr2 0
Rp2 pr2 0 50
Ru2 u2 0 50
Fr2 u2 0 Vsr2 -1
Fu2 u2 0 Vsp2 -1
Ry2 y2 0 1
Gy2 p2 0 y2 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 1.97117285923945
Cx1 x1 xm1 3.07524180660873e-13
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -2.02971788753589
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -0.820391907541706
Cx2 x2 xm2 3.07524180660873e-13
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 1.66516412952709
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 0.370109051834733
Cx3 x3 xm3 6.23727987668804e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -3.29809260983475
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -0.829701297966439
Cx4 x4 xm4 6.23727987668804e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 2.73643171919341
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 2.94812244023603
Cx5 x5 xm5 1.68334113126759e-13
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -1.11219753585198
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -1.39837053340169
Cx6 x6 xm6 1.68334113126759e-13
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 1.55526426145738
Rx7 x7 0 1
Cx7 x7 0 4.45299357322097e-13
Gx7_1 x7 0 u1 0 -2.10997268532332
Rx8 x8 0 1
Cx8 x8 0 3.15154927003678e-12
Gx8_1 x8 0 u1 0 -0.0274521589136151
Rx9 x9 0 1
Cx9 x9 0 1.40481832449782e-11
Gx9_1 x9 0 u1 0 -0.0111541281294792
Rx10 x10 0 1
Fxc10_11 x10 0 Vx11 2.61688157948964
Cx10 x10 xm10 3.07524180660873e-13
Vx10 xm10 0 0
Gx10_2 x10 0 u2 0 -2.04869967256455
Rx11 x11 0 1
Fxc11_10 x11 0 Vx10 -0.617962339129336
Cx11 x11 xm11 3.07524180660873e-13
Vx11 xm11 0 0
Gx11_2 x11 0 u2 0 1.2660192418315
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 0.317692735724175
Cx12 x12 xm12 6.23727987668804e-13
Vx12 xm12 0 0
Gx12_2 x12 0 u2 0 -2.81882130051318
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -0.966594215622912
Cx13 x13 xm13 6.23727987668804e-13
Vx13 xm13 0 0
Gx13_2 x13 0 u2 0 2.7246563639507
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 2.93904995546655
Cx14 x14 xm14 1.68334113126759e-13
Vx14 xm14 0 0
Gx14_2 x14 0 u2 0 -1.11495868903734
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -1.40268713079152
Cx15 x15 xm15 1.68334113126759e-13
Vx15 xm15 0 0
Gx15_2 x15 0 u2 0 1.56393820447686
Rx16 x16 0 1
Cx16 x16 0 4.45299357322097e-13
Gx16_2 x16 0 u2 0 -2.63544354717997
Rx17 x17 0 1
Cx17 x17 0 3.15154927003678e-12
Gx17_2 x17 0 u2 0 -0.0272117440038125
Rx18 x18 0 1
Cx18 x18 0 1.40481832449782e-11
Gx18_2 x18 0 u2 0 -0.0107050957148337
Gyc1_1 y1 0 x1 0 0.197077515897355
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 -0.0896393631148316
Gyc1_5 y1 0 x5 0 -0.243334574601374
Gyc1_6 y1 0 x6 0 -0.0555692141281726
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -0.0946854652007274
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 0.726965964037853
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 1
Gyc1_16 y1 0 x16 0 -0.34798965998787
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -0.711867320699658
Gyc2_1 y2 0 x1 0 1
Gyc2_2 y2 0 x2 0 -0.764870767998925
Gyc2_3 y2 0 x3 0 0.612097406604057
Gyc2_4 y2 0 x4 0 1
Gyc2_5 y2 0 x5 0 -1
Gyc2_6 y2 0 x6 0 1
Gyc2_7 y2 0 x7 0 -0.414558672372795
Gyc2_8 y2 0 x8 0 -1
Gyc2_9 y2 0 x9 0 -0.689973873640247
Gyc2_10 y2 0 x10 0 0.397249714170045
Gyc2_11 y2 0 x11 0 0.828935882572111
Gyc2_12 y2 0 x12 0 1
Gyc2_13 y2 0 x13 0 -0.168682286584248
Gyc2_14 y2 0 x14 0 -0.184995428695174
Gyc2_15 y2 0 x15 0 0.141337739811527
Gyc2_16 y2 0 x16 0 -1
Gyc2_17 y2 0 x17 0 0.0651537249882321
Gyc2_18 y2 0 x18 0 1
.ENDS
