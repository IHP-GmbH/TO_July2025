** sch_path: /ALL/Xschem/LC_VCO/VCO_LC_core.sch
.subckt VCO_LC_core out_n out_p VDD VSS c2 c1 v_gain
*.PININFO VSS:B VDD:B c1:B c2:B out_p:B out_n:B v_gain:B
x2 v_gain c1 c2 c2 c1 VSS dual_inv nw=3e-05 nl=1.3e-07 pw=9e-05 pl=1.3e-07
C2 VSS v_gain cap_cmim w=28e-6 l=18e-6
x1 VDD out_p out_n c1 c2 VSS dual_inv nw=3e-05 nl=1.3e-07 pw=9e-05 pl=1.3e-07
C1 VSS VDD cap_cmim w=28e-6 l=16e-6
**** begin user architecture code




**** end user architecture code
.ends

* expanding   symbol:  /ALL/Xschem/LC_VCO/dual_inv.sym # of pins=6
** sym_path: /ALL/Xschem/LC_VCO/dual_inv.sym
** sch_path: /ALL/Xschem/LC_VCO/dual_inv.sch
.subckt dual_inv VDD out_p out_n in_n in_p VSS  symname=diffamp nw=1u nl=1u pw=2u pl=1u
*.PININFO out_p:B out_n:B in_p:B in_n:B VSS:B VDD:B
**** begin user architecture code


**** end user architecture code
M31 out_p in_n VSS VSS sg13_lv_nmos w={nw} l={nl} m=1 ng=1
M32 out_p in_n VDD VDD sg13_lv_pmos w={pw} l={pl} m=1 ng=1
M49 out_n in_p VSS VSS sg13_lv_nmos w={nw} l={nl} m=1 ng=1
M50 out_n in_p VDD VDD sg13_lv_pmos w={pw} l={pl} m=1 ng=1
.ends

