** sch_path: /ALL/Xschem/LC_VCO/measuremenst_and_test_of_idas/VCO_LC__TB_05_ac_lv_nmosSW.sch
**.subckt VCO_LC__TB_05_ac_lv_nmosSW
VDD VDD GND 1.4
VSS GND VSS 0
Vx6 net2 VSS 0 ac 1 0
C6 VSS net1 1p
L27 net85 net1 2.2n
R1 net85 VSS 3.5
Vx5 net1 VSS 0 ac 1 0
C7 VSS net2 1.2p
L32 net86 net2 2.2n
R3 net86 VSS 3.5
VDD1 0 GND 0
VCO VCO GND .7 pulse(0 2 1n 100n 100n 100n 1)
Vddd1 VCO net3 0
L10 P5 net4 2.2n
R4 net4 N5 3.5
XC1 P5 N5 cap_cmim w=10.0e-6 l=33.0e-6
XC4 P5 N5 cap_cmim w=10.0e-6 l=16.0e-6
XC5 P5 N5 cap_cmim w=10.0e-6 l=8.0e-6
XC8 P5 N5 cap_cmim w=10.0e-6 l=4.0e-6
R7 net5 N5 7.5
C3 net6 net5 120f
C9 net7 net6 120f
R8 P5 net7 7.5
R5 net6 net3 10k
I2 N5 P5 0 ac 1 0
Vddd8 VCO net8 0
L21 P15 net9 2.2n
R14 net9 N15 3.5
XC16 P15 N15 cap_cmim w=10.0e-6 l=16.0e-6
XC17 P15 N15 cap_cmim w=10.0e-6 l=8.0e-6
XC18 P15 N15 cap_cmim w=10.0e-6 l=4.0e-6
R15 net10 N15 7.5
C19 net11 net10 120f
C20 net12 net11 120f
R16 P15 net12 7.5
R17 net11 net8 10k
I3 N15 P15 0 ac 1 0
Vddd11 VCO net13 0
L35 P25 net14 2.2n
R19 net14 N25 3.5
R20 net15 N25 7.5
C25 net16 net15 120f
C26 net17 net16 120f
R22 P25 net17 7.5
R23 net16 net13 10k
I4 N25 P25 0 ac 1 0
XM31 NMOSr1 net18 VSS VSS sg13_lv_nmos w={nsw2} l=.13u ng=1
I5 NMOSr1 VSS 0 ac 1 0
VDD2 net18 VSS 2
XM1 NMOSrO net19 VSS VSS sg13_lv_nmos w={nsw2} l=.13u ng=1
I6 NMOSrO VSS 0 ac 1 0
VDD3 net19 VSS 0
R6 VCO N5 111k
R9 P5 VCO 111k
R10 VCO N15 111k
R11 P15 VCO 111k
R12 VCO N25 111k
R34 P25 VCO 111k
L55 P5s3 net20 2.2n
R69 net20 N5s3 3.5
XC59 net25 net21 cap_cmim w=10.0e-6 l=32.0e-6
R70 net22 N5s3 7.5
C63 net23 net22 120f
C64 net24 net23 120f
R71 P5s3 net24 7.5
R72 net23 VCO 10k
I11 N5s3 P5s3 0 ac 1 0
XM43 net21 net28 N5s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
XM44 net25 net27 P5s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
VDD9 net26 VSS 1.8
R73 VCO N5s3 111k
R74 P5s3 VCO 111k
XC65 net27 P5s3 cap_cmim w=20.0e-6 l=20.0e-6
R75 net26 net27 11k
XC69 net28 N5s3 cap_cmim w=20.0e-6 l=20.0e-6
R79 net28 net26 11k
XM47 VSS net29 VSS VSS sg13_lv_nmos w={nsw2} l=.13u ng=1
VDD11 net29 VSS 0 ac 1 0
XC73 net31 net30 cap_cmim w=10.0e-6 l=16.0e-6
XM88 net30 net33 N5s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XM89 net31 net32 P5s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XC74 net32 P5s3 cap_cmim w=20.0e-6 l=10.0e-6
R116 net26 net32 11k
XC75 net33 N5s3 cap_cmim w=20.0e-6 l=10.0e-6
R117 net33 net26 11k
XC2 net35 net34 cap_cmim w=10.0e-6 l=8.0e-6
XM2 net34 net37 N5s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XM3 net35 net36 P5s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XC10 net36 P5s3 cap_cmim w=20.0e-6 l=5.0e-6
R24 net26 net36 11k
XC11 net37 N5s3 cap_cmim w=20.0e-6 l=5.0e-6
R25 net37 net26 11k
XC12 net39 net38 cap_cmim w=10.0e-6 l=4.0e-6
XM4 net38 net41 N5s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XM5 net39 net40 P5s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XC13 net40 P5s3 cap_cmim w=20.0e-6 l=2.5e-6
R26 net26 net40 11k
XC14 net41 N5s3 cap_cmim w=20.0e-6 l=2.5e-6
R27 net41 net26 11k
L12 P15s3 net42 2.2n
R29 net42 N15s3 3.5
XC27 net47 net43 cap_cmim w=10.0e-6 l=32.0e-6
R30 net44 N15s3 7.5
C28 net45 net44 120f
C29 net46 net45 120f
R31 P15s3 net46 7.5
R32 net45 VCO 10k
I1 N15s3 P15s3 0 ac 1 0
XM6 net43 net50 N15s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
XM7 net47 net49 P15s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
VDD4 net48 VSS 1.8
R33 VCO N15s3 111k
R35 P15s3 VCO 111k
XC30 net49 P15s3 cap_cmim w=20.0e-6 l=20.0e-6
R36 VSS net49 11k
XC31 net50 N15s3 cap_cmim w=20.0e-6 l=20.0e-6
R37 net50 VSS 11k
XC32 net52 net51 cap_cmim w=10.0e-6 l=16.0e-6
XM8 net51 net54 N15s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XM9 net52 net53 P15s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XC33 net53 P15s3 cap_cmim w=20.0e-6 l=10.0e-6
R38 net48 net53 11k
XC34 net54 N15s3 cap_cmim w=20.0e-6 l=10.0e-6
R39 net54 net48 11k
XC35 net56 net55 cap_cmim w=10.0e-6 l=8.0e-6
XM10 net55 net58 N15s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XM11 net56 net57 P15s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XC36 net57 P15s3 cap_cmim w=20.0e-6 l=5.0e-6
R40 net48 net57 11k
XC37 net58 N15s3 cap_cmim w=20.0e-6 l=5.0e-6
R41 net58 net48 11k
XC38 net60 net59 cap_cmim w=10.0e-6 l=4.0e-6
XM12 net59 net62 N15s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XM13 net60 net61 P15s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XC39 net61 P15s3 cap_cmim w=20.0e-6 l=2.5e-6
R42 net48 net61 11k
XC40 net62 N15s3 cap_cmim w=20.0e-6 l=2.5e-6
R43 net62 net48 11k
L23 P25s3 net63 2.2n
R45 net63 N25s3 3.5
XC41 net68 net64 cap_cmim w=10.0e-6 l=32.0e-6
R46 net65 N25s3 7.5
C42 net66 net65 120f
C43 net67 net66 120f
R47 P25s3 net67 7.5
R48 net66 VCO 10k
I7 N25s3 P25s3 0 ac 1 0
XM14 net64 net71 N25s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
XM15 net68 net70 P25s3 VSS sg13_lv_nmos w=480u l=.13u ng=1
VDD5 net69 VSS 0
R49 VCO N25s3 111k
R50 P25s3 VCO 111k
XC44 net70 P25s3 cap_cmim w=20.0e-6 l=20.0e-6
R51 net69 net70 11k
XC45 net71 N25s3 cap_cmim w=20.0e-6 l=20.0e-6
R52 net71 net69 11k
XC46 net73 net72 cap_cmim w=10.0e-6 l=16.0e-6
XM16 net72 net75 N25s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XM17 net73 net74 P25s3 VSS sg13_lv_nmos w=240u l=.13u ng=1
XC47 net74 P25s3 cap_cmim w=20.0e-6 l=10.0e-6
R53 net69 net74 11k
XC48 net75 N25s3 cap_cmim w=20.0e-6 l=10.0e-6
R54 net75 net69 11k
XC49 net77 net76 cap_cmim w=10.0e-6 l=8.0e-6
XM18 net76 net79 N25s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XM19 net77 net78 P25s3 VSS sg13_lv_nmos w=120u l=.13u ng=1
XC50 net78 P25s3 cap_cmim w=20.0e-6 l=5.0e-6
R55 net69 net78 11k
XC51 net79 N25s3 cap_cmim w=20.0e-6 l=5.0e-6
R56 net79 net69 11k
XC52 net81 net80 cap_cmim w=10.0e-6 l=4.0e-6
XM20 net80 net83 N25s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XM21 net81 net82 P25s3 VSS sg13_lv_nmos w=250u l=.13u ng=1
XC53 net82 P25s3 cap_cmim w=20.0e-6 l=2.5e-6
R57 net69 net82 11k
XC54 net83 N25s3 cap_cmim w=20.0e-6 l=2.5e-6
R58 net83 net69 11k
XD1 VDD net84 VSS diodevdd_2kv
XD2 VDD net84 VSS diodevss_2kv
VDD6 net84 VSS 0.7 ac 1 0
**** begin user architecture code







* schematic: VCO_LC__TB_05_ac_lv_nmosSW
* dir:       LC_VCO/measuremenst_and_test_of_idas
* test:      LC_VCO/measuremenst_and_test_of_idas/OTA33_BiAS.sym

* mos_corner:
* mos_corner:






.option temp=27


.inc /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/sg13g2_bondpad.lib
.inc /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/sg13g2_esd.lib
.inc /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/diodes.lib

.lib /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/cornerRES.lib     res_typ
.lib /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/cornerCAP.lib     cap_typ

.lib /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/cornerMOShv.lib   mos_tt
.lib /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/cornerMOSlv.lib   mos_tt
.lib /home/ich/share/pdk/dev/IHP-Open-PDK/ihp-sg13g2/libs.tech/xyce/models/cornerHBT.lib     hbt_typ

.param nw=5e-6
.param nl=.13e-6
.param pw=10e-6
.param pl=.13e-6
.param iset=0

.param nsw2=500u
.param nsw1=100u
.param nsw=50u


*.step vco 0 1.8 .1
.ac dec 111 10e6 101e9
.print ac format=raw v(*) i(*)




**** end user architecture code
**.ends
.GLOBAL GND
.end
